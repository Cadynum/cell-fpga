../nexys3/cell1d/ipcore_dir/clockgen.vhd